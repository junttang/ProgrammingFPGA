`timescale 1ns / 1ps

module inv(
    input a,
    output y
    );
    
    assign y=~a;
endmodule
